-- vou dar um commit antes de iniciar o top-level
